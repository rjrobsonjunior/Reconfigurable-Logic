lpm_counter_ex_inst : lpm_counter_ex PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
