-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Tue Sep 16 17:43:27 2025

FSM_LineFollower FSM_LineFollower_inst
(
	.clock(clock_sig) ,	// input  clock_sig
	.reset(reset_sig) ,	// input  reset_sig
	.LeftSensor(LeftSensor_sig) ,	// input  LeftSensor_sig
	.RightSensor(RightSensor_sig) ,	// input  RightSensor_sig
	.Enable(Enable_sig) ,	// input  Enable_sig
	.Losting(Losting_sig) ,	// input  Losting_sig
	.MotorSpeedLeft(MotorSpeedLeft_sig) ,	// output  MotorSpeedLeft_sig
	.MotorSpeedRight(MotorSpeedRight_sig) ,	// output  MotorSpeedRight_sig
	.Looking(Looking_sig) ,	// output  Looking_sig
	.EnableMotorLeft(EnableMotorLeft_sig) ,	// output  EnableMotorLeft_sig
	.EnableMotorRight(EnableMotorRight_sig) 	// output  EnableMotorRight_sig
);

