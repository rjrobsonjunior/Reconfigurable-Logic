CounterwAclr_inst : CounterwAclr PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
