counter25pins_inst : counter25pins PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
