Mem256sword16bits_inst : Mem256sword16bits PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
