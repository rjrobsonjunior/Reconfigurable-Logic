SQRT32_inst : SQRT32 PORT MAP (
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
