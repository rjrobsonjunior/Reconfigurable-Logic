-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Tue Sep 09 17:06:48 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachineMotor IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        Enable : IN STD_LOGIC := '0';
        Sentido : IN STD_LOGIC := '0';
        Saida1 : OUT STD_LOGIC;
        Saida2 : OUT STD_LOGIC
    );
END StateMachineMotor;

ARCHITECTURE BEHAVIOR OF StateMachineMotor IS
    TYPE type_fstate IS (S1,S2,S3,S0);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_Saida1 : STD_LOGIC := '0';
    SIGNAL reg_Saida2 : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate,reg_Saida1,reg_Saida2)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
            Saida1 <= reg_Saida1;
            Saida2 <= reg_Saida2;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Enable,Sentido)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S0;
            reg_Saida1 <= '0';
            reg_Saida2 <= '0';
        ELSE
            reg_Saida1 <= '0';
            reg_Saida2 <= '0';
            CASE fstate IS
                WHEN S1 =>
                    IF (((Sentido = '1') AND (Enable = '1'))) THEN
                        reg_fstate <= S2;
                    ELSIF (NOT((Enable = '1'))) THEN
                        reg_fstate <= S1;
                    ELSIF ((NOT((Sentido = '1')) AND (Enable = '1'))) THEN
                        reg_fstate <= S0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S1;
                    END IF;

                    reg_Saida2 <= '0';

                    reg_Saida1 <= '1';
                WHEN S2 =>
                    IF (((Sentido = '1') AND (Enable = '1'))) THEN
                        reg_fstate <= S3;
                    ELSIF (NOT((Enable = '1'))) THEN
                        reg_fstate <= S2;
                    ELSIF ((NOT((Sentido = '1')) AND (Enable = '1'))) THEN
                        reg_fstate <= S1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S2;
                    END IF;

                    reg_Saida2 <= '0';

                    reg_Saida1 <= '0';
                WHEN S3 =>
                    IF (((Sentido = '1') AND (Enable = '1'))) THEN
                        reg_fstate <= S0;
                    ELSIF ((NOT((Sentido = '1')) AND (Enable = '1'))) THEN
                        reg_fstate <= S2;
                    ELSIF (NOT((Enable = '1'))) THEN
                        reg_fstate <= S3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S3;
                    END IF;

                    reg_Saida2 <= '1';

                    reg_Saida1 <= '0';
                WHEN S0 =>
                    IF (((Sentido = '1') AND (Enable = '1'))) THEN
                        reg_fstate <= S1;
                    ELSIF (NOT((Enable = '1'))) THEN
                        reg_fstate <= S0;
                    ELSIF ((NOT((Sentido = '1')) AND (Enable = '1'))) THEN
                        reg_fstate <= S3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    reg_Saida2 <= '1';

                    reg_Saida1 <= '1';
                WHEN OTHERS => 
                    reg_Saida1 <= 'X';
                    reg_Saida2 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
