-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Tue Sep 16 17:42:37 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FSM_LineFollower IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        LeftSensor : IN STD_LOGIC := '0';
        RightSensor : IN STD_LOGIC := '0';
        Enable : IN STD_LOGIC := '0';
        Losting : IN STD_LOGIC := '0';
        MotorSpeedLeft : OUT STD_LOGIC;
        MotorSpeedRight : OUT STD_LOGIC;
        Looking : OUT STD_LOGIC;
        EnableMotorLeft : OUT STD_LOGIC;
        EnableMotorRight : OUT STD_LOGIC
    );
END FSM_LineFollower;

ARCHITECTURE BEHAVIOR OF FSM_LineFollower IS
    TYPE type_fstate IS (Idle,FullSpeed,TurnLeft,TurnRight,SeekLeft,SeekRight,Lost);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_MotorSpeedLeft : STD_LOGIC := '0';
    SIGNAL reg_MotorSpeedRight : STD_LOGIC := '0';
    SIGNAL reg_Looking : STD_LOGIC := '0';
    SIGNAL reg_EnableMotorLeft : STD_LOGIC := '0';
    SIGNAL reg_EnableMotorRight : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate,reg_MotorSpeedLeft,reg_MotorSpeedRight,reg_Looking,reg_EnableMotorLeft)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
            MotorSpeedLeft <= reg_MotorSpeedLeft;
            MotorSpeedRight <= reg_MotorSpeedRight;
            Looking <= reg_Looking;
            EnableMotorLeft <= reg_EnableMotorLeft;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,LeftSensor,RightSensor,Enable,Losting,reg_EnableMotorRight)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Idle;
            reg_MotorSpeedLeft <= '0';
            reg_MotorSpeedRight <= '0';
            reg_Looking <= '0';
            reg_EnableMotorLeft <= '0';
            reg_EnableMotorRight <= '0';
            EnableMotorRight <= '0';
        ELSE
            reg_MotorSpeedLeft <= '0';
            reg_MotorSpeedRight <= '0';
            reg_Looking <= '0';
            reg_EnableMotorLeft <= '0';
            reg_EnableMotorRight <= '0';
            EnableMotorRight <= '0';
            CASE fstate IS
                WHEN Idle =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    ELSIF (((Enable = '1') AND (Losting = '1'))) THEN
                        reg_fstate <= Lost;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= SeekRight;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Idle;
                    END IF;

                    reg_MotorSpeedRight <= '0';

                    reg_Looking <= '0';

                    reg_EnableMotorLeft <= '0';
                    reg_EnableMotorLeft <= '0';

                    reg_MotorSpeedLeft <= '0';

                    reg_EnableMotorRight <= '0';
                WHEN FullSpeed =>
                    IF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= SeekRight;
                    ELSIF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= FullSpeed;
                    END IF;

                    reg_MotorSpeedRight <= '1';

                    reg_Looking <= '0';

                    reg_EnableMotorLeft <= '1';

                    reg_MotorSpeedLeft <= '1';

                    reg_EnableMotorRight <= '1';
                WHEN TurnLeft =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= SeekLeft;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= TurnLeft;
                    END IF;

                    reg_MotorSpeedRight <= '0';

                    reg_Looking <= '0';

                    reg_EnableMotorLeft <= '1';

                    reg_MotorSpeedLeft <= '1';

                    reg_EnableMotorRight <= '1';
                WHEN TurnRight =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= SeekRight;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= TurnRight;
                    END IF;

                    reg_MotorSpeedRight <= '1';

                    reg_Looking <= '0';

                    reg_EnableMotorLeft <= '1';

                    reg_MotorSpeedLeft <= '0';

                    reg_EnableMotorRight <= '1';
                WHEN SeekLeft =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    ELSIF (((Enable = '1') AND (Losting = '1'))) THEN
                        reg_fstate <= Lost;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SeekLeft;
                    END IF;

                    reg_MotorSpeedRight <= '0';

                    reg_Looking <= '0';

                    reg_EnableMotorLeft <= '1';

                    reg_MotorSpeedLeft <= '1';

                    reg_EnableMotorRight <= '0';
                WHEN SeekRight =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND (RightSensor = '1'))) THEN
                        reg_fstate <= FullSpeed;
                    ELSIF (((Enable = '1') AND (Losting = '1'))) THEN
                        reg_fstate <= Lost;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND NOT((LeftSensor = '1'))) AND (RightSensor = '1'))) THEN
                        reg_fstate <= TurnLeft;
                    ELSIF (((((Enable = '1') AND NOT((Losting = '1'))) AND (LeftSensor = '1')) AND NOT((RightSensor = '1')))) THEN
                        reg_fstate <= TurnRight;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SeekRight;
                    END IF;

                    reg_MotorSpeedRight <= '1';

                    reg_Looking <= '1';

                    reg_EnableMotorLeft <= '0';

                    reg_MotorSpeedLeft <= '0';

                    reg_EnableMotorRight <= '1';
                WHEN Lost =>
                    IF (NOT((Enable = '1'))) THEN
                        reg_fstate <= Idle;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Lost;
                    END IF;

                    reg_MotorSpeedRight <= '0';

                    reg_Looking <= '0';

                    reg_MotorSpeedLeft <= '0';

                    reg_EnableMotorRight <= '0';
                WHEN OTHERS => 
                    reg_MotorSpeedLeft <= 'X';
                    reg_MotorSpeedRight <= 'X';
                    reg_Looking <= 'X';
                    reg_EnableMotorLeft <= 'X';
                    reg_EnableMotorRight <= 'X';
                    report "Reach undefined state";
            END CASE;
            EnableMotorRight <= reg_EnableMotorRight;
        END IF;
    END PROCESS;
END BEHAVIOR;
