Counter16_inst : Counter16 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
