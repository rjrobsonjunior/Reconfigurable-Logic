Counter10s_inst : Counter10s PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
